`define IF_TO_ID_WD 33
`define ID_TO_EX_WD 149
`define EX_TO_MEM_WD 76
`define MEM_TO_WB_WD 271
`define BR_WD 33
`define DATA_SRAM_WD 69
`define WB_TO_RF_WD 38

`define StallBus 6
`define NoStop 1'b0
`define Stop 1'b1