`include "defines.vh"
module WB(
    input wire clk,
    input wire rst
);
    
endmodule