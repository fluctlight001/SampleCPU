`include "lib/defines.vh"
module CTRL(
    input wire rst,
    input wire stallreq_from
);

endmodule