`include "defines.vh"
module MEM(
    input wire clk,
    input wire rst
);
    
endmodule